library verilog;
use verilog.vl_types.all;
entity Diretorio is
    port(
        Clock           : in     vl_logic
    );
end Diretorio;
