library verilog;
use verilog.vl_types.all;
entity Processador2 is
    port(
        Clock           : in     vl_logic;
        AddressTest     : in     vl_logic_vector(3 downto 0);
        WriteOrRead     : in     vl_logic_vector(2 downto 0);
        Processor       : in     vl_logic_vector(2 downto 0);
        DataTest        : in     vl_logic_vector(3 downto 0);
        HitOrMissP2     : out    vl_logic_vector(1 downto 0);
        HitOrMissP1     : in     vl_logic_vector(1 downto 0);
        WriteBack       : out    vl_logic_vector(1 downto 0)
    );
end Processador2;
